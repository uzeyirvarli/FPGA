----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:06:07 04/15/2020 
-- Design Name: 
-- Module Name:    FSM_Moore_Code2 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity FSM_Moore_Code2 is
    Port ( w : in  STD_LOGIC;
           clock  : in  STD_LOGIC;
           Resetn : in  STD_LOGIC;
           z : out  STD_LOGIC);
end FSM_Moore_Code2;

architecture Behavioral of FSM_Moore_Code2 is

begin


end Behavioral;

